*** SPICE deck for cell regulation_circuit{sch} from library Lab_06
*** Created on Thu Nov 06, 2025 19:56:33
*** Last revised on Thu Nov 06, 2025 20:23:02
*** Written on Thu Nov 06, 2025 23:06:12 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: regulation_circuit{sch}
Mnmos@0 net@21 net@9 gnd gnd N_50n L=0.3U W=3U
Mnmos@1 net@24 net@21 gnd gnd N_50n L=0.3U W=3U
Mnmos@2 En net@24 gnd gnd N_50n L=0.3U W=3U
Mpmos@0 net@21 gnd vdd vdd P_50n L=12U W=6U
Mpmos@1 net@21 net@24 vdd vdd P_50n L=12U W=6U
Mpmos@2 net@24 net@21 vdd vdd P_50n L=0.3U W=6U
Mpmos@3 En net@24 vdd vdd P_50n L=0.3U W=6U
Rres@0 vdd net@9 20MEG
Rres@1 net@9 Vout 3MEG

* Spice Code nodes in cell cell 'regulation_circuit{sch}'
vdd vdd 0 DC 1V
vout vout 0 SIN(1.5 1.5 50)
.tran 0 1
.include cmosedu_models.txt
.END
