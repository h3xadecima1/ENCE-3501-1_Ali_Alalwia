*** SPICE deck for cell XOR_Gate_SIM_2{sch} from library Lab_05
*** Created on Fri Oct 24, 2025 19:24:13
*** Last revised on Fri Oct 24, 2025 19:29:55
*** Written on Fri Oct 24, 2025 19:30:00 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Lab_05__XOR_Gate FROM CELL XOR_Gate{sch}
.SUBCKT Lab_05__XOR_Gate A AxorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@63 B gnd gnd NMOS L=0.6U W=1.8U
Mnmos@1 net@64 net@120 gnd gnd NMOS L=0.6U W=1.8U
Mnmos@2 AxorB A net@63 gnd NMOS L=0.6U W=1.8U
Mnmos@3 AxorB net@144 net@64 gnd NMOS L=0.6U W=1.8U
Mnmos@4 net@120 B gnd gnd NMOS L=0.6U W=1.8U
Mnmos@5 net@144 A gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd A net@46 vdd PMOS L=0.6U W=1.8U
Mpmos@1 vdd B net@46 vdd PMOS L=0.6U W=1.8U
Mpmos@2 net@46 net@144 AxorB vdd PMOS L=0.6U W=1.8U
Mpmos@3 net@46 net@120 AxorB vdd PMOS L=0.6U W=1.8U
Mpmos@4 vdd B net@120 vdd PMOS L=0.6U W=1.8U
Mpmos@5 vdd A net@144 vdd PMOS L=0.6U W=1.8U
.ENDS Lab_05__XOR_Gate

.global gnd vdd

*** TOP LEVEL CELL: XOR_Gate_SIM_2{sch}
XXOR_Gate@0 d_in exor_out vdd Lab_05__XOR_Gate

* Spice Code nodes in cell cell 'XOR_Gate_SIM_2{sch}'
vdd vdd 0 dc 5
vin d_in 0 pulse(0v 5v 10n 1n 1n 40n 42n)
.tran 0 40n
.include C5_models.txt
.END
