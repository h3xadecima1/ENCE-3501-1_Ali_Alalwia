*** SPICE deck for cell NOT_Gate_SIM{sch} from library Lab_05
*** Created on Fri Oct 24, 2025 16:26:28
*** Last revised on Fri Oct 24, 2025 16:28:16
*** Written on Fri Oct 24, 2025 16:28:21 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Lab_05__NOT_Gate FROM CELL NOT_Gate{sch}
.SUBCKT Lab_05__NOT_Gate In Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out In gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd In Out vdd PMOS L=0.6U W=1.8U
.ENDS Lab_05__NOT_Gate

.global gnd vdd

*** TOP LEVEL CELL: NOT_Gate_SIM{sch}
XNOT_Gate@0 d_in not_d_out Lab_05__NOT_Gate

* Spice Code nodes in cell cell 'NOT_Gate_SIM{sch}'
vdd vdd 0 dc 5
vin d_in 0 pulse(0v 5v 10n 1n 1n 40n 42n)
.tran 0 40n
.include C5_models.txt
.END
